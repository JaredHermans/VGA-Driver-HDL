//The purpose of this module is to modify the input HSync and VSync signals to
//include some time for what is called the Front and Back porch. The front and 
//back porch of a VGA interfase used to have more meaning when a monitor
//actually used a Cathode Ray Tube (CRT) to draw an image on the screen. New 
//standards like DVI and HDMI which are meant for digital signals have
//removed this notion of the front and back porches. Remember that VGA is an analog
//interface.
//This module is designed for 640 x 480 with a 25 MHz input clock

module VGA_Sync_Porch #(
    parameter                       VIDEO_WIDTH = 3,
    parameter                       TOTAL_COLS  = 3,
    parameter                       TOTAL_ROWS  = 3,
    parameter                       ACTIVE_COLS = 3,
    parameter                       ACTIVE_ROWS = 3
)
(
    input                           i_Clk,
    input                           i_HSync,
    input                           i_VSync,
    input [VIDEO_WIDTH - 1:0]       i_Red_Video,
    input [VIDEO_WIDTH - 1:0]       i_Grn_Video,
    input [VIDEO_WIDTH - 1:0]       i_Blu_Video,
    output reg                      o_HSync,
    output reg                      o_VSync,
    output reg [VIDEO_WIDTH - 1:0]  o_Red_Video,
    output reg [VIDEO_WIDTH - 1:0]  o_Grn_Video,
    output reg [VIDEO_WIDTH - 1:0]  o_Blu_Video 
);
    parameter c_FRONT_PORCH_HORZ    = 21;
    parameter c_BACK_PORCH_HORZ     = 48;
    parameter c_FRONT_PORCH_VERT    = 8;
    parameter c_BACK_PORCH_VERT     = 36;

    wire w_HSync;
    wire w_VSync;

    wire [9:0] w_Col_Count;
    wire [9:0] w_Row_Count;

    reg [VIDEO_WIDTH - 1:0] r_Red_Video = 0;
    reg [VIDEO_WIDTH - 1:0] r_Grn_Video = 0;
    reg [VIDEO_WIDTH - 1:0] r_Blu_Video = 0;

    Sync_To_Count #(
        .TOTAL_COLS     (TOTAL_COLS),
        .TOTAL_ROWS     (TOTAL_ROWS)
    )
    UUT (
        .i_Clk          (i_Clk),
        .i_HSync        (i_HSync),
        .i_VSync        (i_VSync),
        .o_HSync        (w_HSync),
        .o_VSync        (w_VSync),
        .o_Col_Count    (w_Col_Count),
        .o_Row_Count    (w_Row_Count)
    );

    //Purpose: Modifies the HSync and VSync signals to include Front/Back porch
    always @ (posedge i_Clk) begin
        if ((w_Col_Count < c_FRONT_PORCH_HORZ + ACTIVE_COLS) || (w_Col_Count > TOTAL_COLS - c_BACK_PORCH_HORZ - 1))
            o_HSync <= 1'b1;
        else
            o_HSync <= w_HSync;

        if ((w_Row_Count < c_FRONT_PORCH_VERT + ACTIVE_ROWS) || (w_Row_Count > TOTAL_ROWS - c_BACK_PORCH_VERT - 1))
            o_VSync <=  1'b1;
        else 
            o_VSync <= w_VSync; 
    end

    //Purpose: Align input video to modified Sync Pulses.
    //Adds in 2 Clock Cycles of Deley
    always @ (posedge i_Clk) begin
        r_Red_Video <= i_Red_Video;
        r_Grn_Video <= i_Grn_Video;
        r_Blu_Video <= i_Blu_Video;

        o_Red_Video <= r_Red_Video;
        o_Grn_Video <= r_Grn_Video;
        o_Blu_Video <= r_Blu_Video;
    end

endmodule